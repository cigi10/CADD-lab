`timescale 1ns / 1ps

module mux_2_1
    (
    input wire d0,     
    input wire d1,     
    input wire s,      
    output wire y      
);
    assign y = s ? d1 : d0;
endmodule
